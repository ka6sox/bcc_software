`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:07:30 06/12/2013 
// Design Name: 
// Module Name:    gpmc_sram 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module gpmc_sram(
		input			 GPMC_CLK,
		inout [15:0] GPMC_AD,
		input	       GPMC_CS,
		input        GPMC_ADV,
		input			 GPMC_OE,
		input			 GPMC_WE,
		input			 GPMC_BE0,
		input			 GPMC_BE1,
		input			 GPMC_WP,
		input			 GPMC_DIR
);




endmodule
